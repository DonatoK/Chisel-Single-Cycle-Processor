module control_unit( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input        io_clock, // @[:@6.4]
  input        io_reset, // @[:@6.4]
  input  [6:0] io_opcode, // @[:@6.4]
  output       io_branch_op, // @[:@6.4]
  output       io_memRead, // @[:@6.4]
  output       io_memtoReg, // @[:@6.4]
  output [2:0] io_ALUOp, // @[:@6.4]
  output [1:0] io_next_PC_sel, // @[:@6.4]
  output [1:0] io_operand_A_sel, // @[:@6.4]
  output       io_operand_B_sel, // @[:@6.4]
  output [1:0] io_extend_sel, // @[:@6.4]
  output       io_memWrite, // @[:@6.4]
  output       io_regWrite // @[:@6.4]
);
  wire  _T_31; // @[control_unit.scala 43:20:@8.4]
  wire  _T_32; // @[control_unit.scala 43:46:@9.4]
  wire  _T_33; // @[control_unit.scala 43:32:@10.4]
  wire  _T_34; // @[control_unit.scala 43:72:@11.4]
  wire  _T_35; // @[control_unit.scala 43:58:@12.4]
  wire  _T_36; // @[control_unit.scala 44:23:@13.4]
  wire  _T_37; // @[control_unit.scala 44:9:@14.4]
  wire  _T_38; // @[control_unit.scala 44:47:@15.4]
  wire  _T_39; // @[control_unit.scala 44:33:@16.4]
  wire  _T_40; // @[control_unit.scala 44:70:@17.4]
  wire  _T_41; // @[control_unit.scala 44:56:@18.4]
  wire  _T_42; // @[control_unit.scala 45:23:@19.4]
  wire  _T_46; // @[control_unit.scala 51:19:@27.4]
  wire  _T_49; // @[control_unit.scala 57:19:@34.4]
  wire  _T_70; // @[control_unit.scala 85:38:@82.14]
  wire  _T_74; // @[control_unit.scala 87:38:@89.16]
  wire [2:0] _GEN_5; // @[control_unit.scala 87:61:@90.16]
  wire [2:0] _GEN_6; // @[control_unit.scala 85:61:@83.14]
  wire [2:0] _GEN_7; // @[control_unit.scala 83:37:@76.12]
  wire [2:0] _GEN_8; // @[control_unit.scala 81:35:@71.10]
  wire [2:0] _GEN_9; // @[control_unit.scala 79:36:@66.8]
  wire [2:0] _GEN_10; // @[control_unit.scala 77:37:@61.6]
  wire [1:0] _GEN_12; // @[control_unit.scala 97:61:@109.8]
  wire [1:0] _GEN_13; // @[control_unit.scala 95:34:@102.6]
  wire  _T_88; // @[control_unit.scala 103:33:@117.4]
  wire  _T_90; // @[control_unit.scala 103:57:@119.4]
  wire  _T_92; // @[control_unit.scala 104:31:@121.4]
  wire  _T_99; // @[control_unit.scala 111:33:@132.4]
  wire [1:0] _GEN_17; // @[control_unit.scala 113:38:@138.6]
  wire [1:0] _GEN_19; // @[control_unit.scala 125:36:@162.8]
  wire [1:0] _GEN_20; // @[control_unit.scala 123:36:@157.6]
  assign _T_31 = io_opcode == 7'h33; // @[control_unit.scala 43:20:@8.4]
  assign _T_32 = io_opcode == 7'h13; // @[control_unit.scala 43:46:@9.4]
  assign _T_33 = _T_31 | _T_32; // @[control_unit.scala 43:32:@10.4]
  assign _T_34 = io_opcode == 7'h3; // @[control_unit.scala 43:72:@11.4]
  assign _T_35 = _T_33 | _T_34; // @[control_unit.scala 43:58:@12.4]
  assign _T_36 = io_opcode == 7'h67; // @[control_unit.scala 44:23:@13.4]
  assign _T_37 = _T_35 | _T_36; // @[control_unit.scala 44:9:@14.4]
  assign _T_38 = io_opcode == 7'h6f; // @[control_unit.scala 44:47:@15.4]
  assign _T_39 = _T_37 | _T_38; // @[control_unit.scala 44:33:@16.4]
  assign _T_40 = io_opcode == 7'h17; // @[control_unit.scala 44:70:@17.4]
  assign _T_41 = _T_39 | _T_40; // @[control_unit.scala 44:56:@18.4]
  assign _T_42 = io_opcode == 7'h37; // @[control_unit.scala 45:23:@19.4]
  assign _T_46 = io_opcode == 7'h23; // @[control_unit.scala 51:19:@27.4]
  assign _T_49 = io_opcode == 7'h63; // @[control_unit.scala 57:19:@34.4]
  assign _T_70 = _T_36 | _T_38; // @[control_unit.scala 85:38:@82.14]
  assign _T_74 = _T_40 | _T_42; // @[control_unit.scala 87:38:@89.16]
  assign _GEN_5 = _T_74 ? 3'h6 : 3'h0; // @[control_unit.scala 87:61:@90.16]
  assign _GEN_6 = _T_70 ? 3'h3 : _GEN_5; // @[control_unit.scala 85:61:@83.14]
  assign _GEN_7 = _T_49 ? 3'h2 : _GEN_6; // @[control_unit.scala 83:37:@76.12]
  assign _GEN_8 = _T_34 ? 3'h4 : _GEN_7; // @[control_unit.scala 81:35:@71.10]
  assign _GEN_9 = _T_46 ? 3'h5 : _GEN_8; // @[control_unit.scala 79:36:@66.8]
  assign _GEN_10 = _T_32 ? 3'h1 : _GEN_9; // @[control_unit.scala 77:37:@61.6]
  assign _GEN_12 = _T_70 ? 2'h2 : 2'h0; // @[control_unit.scala 97:61:@109.8]
  assign _GEN_13 = _T_42 ? 2'h3 : _GEN_12; // @[control_unit.scala 95:34:@102.6]
  assign _T_88 = _T_32 | _T_46; // @[control_unit.scala 103:33:@117.4]
  assign _T_90 = _T_88 | _T_34; // @[control_unit.scala 103:57:@119.4]
  assign _T_92 = _T_90 | _T_40; // @[control_unit.scala 104:31:@121.4]
  assign _T_99 = _T_32 | _T_34; // @[control_unit.scala 111:33:@132.4]
  assign _GEN_17 = _T_46 ? 2'h1 : 2'h2; // @[control_unit.scala 113:38:@138.6]
  assign _GEN_19 = _T_36 ? 2'h3 : 2'h0; // @[control_unit.scala 125:36:@162.8]
  assign _GEN_20 = _T_38 ? 2'h2 : _GEN_19; // @[control_unit.scala 123:36:@157.6]
  assign io_branch_op = io_opcode == 7'h63; // @[control_unit.scala 58:18:@36.6 control_unit.scala 60:18:@39.6]
  assign io_memRead = io_opcode == 7'h3; // @[control_unit.scala 64:16:@43.6 control_unit.scala 66:16:@46.6]
  assign io_memtoReg = io_opcode == 7'h3; // @[control_unit.scala 70:17:@50.6 control_unit.scala 72:17:@53.6]
  assign io_ALUOp = _T_31 ? 3'h0 : _GEN_10; // @[control_unit.scala 76:14:@57.6 control_unit.scala 78:14:@62.8 control_unit.scala 80:14:@67.10 control_unit.scala 82:14:@72.12 control_unit.scala 84:14:@77.14 control_unit.scala 86:14:@84.16 control_unit.scala 88:14:@91.18 control_unit.scala 90:14:@94.18]
  assign io_next_PC_sel = _T_49 ? 2'h1 : _GEN_20; // @[control_unit.scala 122:20:@153.6 control_unit.scala 124:20:@158.8 control_unit.scala 126:20:@163.10 control_unit.scala 128:21:@166.10]
  assign io_operand_A_sel = _T_40 ? 2'h1 : _GEN_13; // @[control_unit.scala 94:22:@98.6 control_unit.scala 96:22:@103.8 control_unit.scala 98:22:@110.10 control_unit.scala 100:22:@113.10]
  assign io_operand_B_sel = _T_92 | _T_42; // @[control_unit.scala 106:22:@125.6 control_unit.scala 108:22:@128.6]
  assign io_extend_sel = _T_99 ? 2'h0 : _GEN_17; // @[control_unit.scala 112:19:@134.6 control_unit.scala 114:19:@139.8 control_unit.scala 116:19:@146.10 control_unit.scala 118:19:@149.10]
  assign io_memWrite = io_opcode == 7'h23; // @[control_unit.scala 52:18:@29.6 control_unit.scala 54:18:@32.6]
  assign io_regWrite = _T_41 | _T_42; // @[control_unit.scala 46:18:@22.6 control_unit.scala 48:18:@25.6]
endmodule
