module register_file( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_clock, // @[:@6.4]
  input         io_reset, // @[:@6.4]
  input         io_wEn, // @[:@6.4]
  input  [31:0] io_write_data, // @[:@6.4]
  input  [4:0]  io_read_sel1, // @[:@6.4]
  input  [4:0]  io_read_sel2, // @[:@6.4]
  input  [4:0]  io_write_sel, // @[:@6.4]
  output [31:0] io_read_data1, // @[:@6.4]
  output [31:0] io_read_data2 // @[:@6.4]
);
  reg [31:0] register_file_block_0; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_0;
  reg [31:0] register_file_block_1; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_1;
  reg [31:0] register_file_block_2; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_2;
  reg [31:0] register_file_block_3; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_3;
  reg [31:0] register_file_block_4; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_4;
  reg [31:0] register_file_block_5; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_5;
  reg [31:0] register_file_block_6; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_6;
  reg [31:0] register_file_block_7; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_7;
  reg [31:0] register_file_block_8; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_8;
  reg [31:0] register_file_block_9; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_9;
  reg [31:0] register_file_block_10; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_10;
  reg [31:0] register_file_block_11; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_11;
  reg [31:0] register_file_block_12; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_12;
  reg [31:0] register_file_block_13; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_13;
  reg [31:0] register_file_block_14; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_14;
  reg [31:0] register_file_block_15; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_15;
  reg [31:0] register_file_block_16; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_16;
  reg [31:0] register_file_block_17; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_17;
  reg [31:0] register_file_block_18; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_18;
  reg [31:0] register_file_block_19; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_19;
  reg [31:0] register_file_block_20; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_20;
  reg [31:0] register_file_block_21; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_21;
  reg [31:0] register_file_block_22; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_22;
  reg [31:0] register_file_block_23; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_23;
  reg [31:0] register_file_block_24; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_24;
  reg [31:0] register_file_block_25; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_25;
  reg [31:0] register_file_block_26; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_26;
  reg [31:0] register_file_block_27; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_27;
  reg [31:0] register_file_block_28; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_28;
  reg [31:0] register_file_block_29; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_29;
  reg [31:0] register_file_block_30; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_30;
  reg [31:0] register_file_block_31; // @[regFile.scala 28:32:@8.4]
  reg [31:0] _RAND_31;
  wire  _T_60; // @[regFile.scala 30:15:@9.4]
  wire  _T_67; // @[regFile.scala 34:43:@18.8]
  wire  _T_68; // @[regFile.scala 34:26:@19.8]
  wire [31:0] _GEN_0; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_1; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_2; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_3; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_4; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_5; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_6; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_7; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_8; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_9; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_10; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_11; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_12; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_13; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_14; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_15; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_16; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_17; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_18; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_19; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_20; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_21; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_22; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_23; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_24; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_25; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_26; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_27; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_28; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_29; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_30; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_31; // @[regFile.scala 35:43:@21.10]
  wire [31:0] _GEN_32; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_33; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_34; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_35; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_36; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_37; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_38; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_39; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_40; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_41; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_42; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_43; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_44; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_45; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_46; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_47; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_48; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_49; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_50; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_51; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_52; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_53; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_54; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_55; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_56; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_57; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_58; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_59; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_60; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_61; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_62; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_63; // @[regFile.scala 34:53:@20.8]
  wire [31:0] _GEN_64; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_65; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_66; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_67; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_68; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_69; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_70; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_71; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_72; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_73; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_74; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_75; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_76; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_77; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_78; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_79; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_80; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_81; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_82; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_83; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_84; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_85; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_86; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_87; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_88; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_89; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_90; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_91; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_92; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_93; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_94; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_95; // @[regFile.scala 31:23:@13.6]
  wire [31:0] _GEN_129; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_130; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_131; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_132; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_133; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_134; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_135; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_136; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_137; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_138; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_139; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_140; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_141; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_142; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_143; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_144; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_145; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_146; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_147; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_148; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_149; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_150; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_151; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_152; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_153; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_154; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_155; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_156; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_157; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_158; // @[regFile.scala 43:17:@28.4]
  wire [31:0] _GEN_161; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_162; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_163; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_164; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_165; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_166; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_167; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_168; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_169; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_170; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_171; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_172; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_173; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_174; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_175; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_176; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_177; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_178; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_179; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_180; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_181; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_182; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_183; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_184; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_185; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_186; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_187; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_188; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_189; // @[regFile.scala 44:17:@29.4]
  wire [31:0] _GEN_190; // @[regFile.scala 44:17:@29.4]
  assign _T_60 = $unsigned(clock); // @[regFile.scala 30:15:@9.4]
  assign _T_67 = io_write_sel != 5'h0; // @[regFile.scala 34:43:@18.8]
  assign _T_68 = io_wEn & _T_67; // @[regFile.scala 34:26:@19.8]
  assign _GEN_0 = 5'h0 == io_write_sel ? io_write_data : register_file_block_0; // @[regFile.scala 35:43:@21.10]
  assign _GEN_1 = 5'h1 == io_write_sel ? io_write_data : register_file_block_1; // @[regFile.scala 35:43:@21.10]
  assign _GEN_2 = 5'h2 == io_write_sel ? io_write_data : register_file_block_2; // @[regFile.scala 35:43:@21.10]
  assign _GEN_3 = 5'h3 == io_write_sel ? io_write_data : register_file_block_3; // @[regFile.scala 35:43:@21.10]
  assign _GEN_4 = 5'h4 == io_write_sel ? io_write_data : register_file_block_4; // @[regFile.scala 35:43:@21.10]
  assign _GEN_5 = 5'h5 == io_write_sel ? io_write_data : register_file_block_5; // @[regFile.scala 35:43:@21.10]
  assign _GEN_6 = 5'h6 == io_write_sel ? io_write_data : register_file_block_6; // @[regFile.scala 35:43:@21.10]
  assign _GEN_7 = 5'h7 == io_write_sel ? io_write_data : register_file_block_7; // @[regFile.scala 35:43:@21.10]
  assign _GEN_8 = 5'h8 == io_write_sel ? io_write_data : register_file_block_8; // @[regFile.scala 35:43:@21.10]
  assign _GEN_9 = 5'h9 == io_write_sel ? io_write_data : register_file_block_9; // @[regFile.scala 35:43:@21.10]
  assign _GEN_10 = 5'ha == io_write_sel ? io_write_data : register_file_block_10; // @[regFile.scala 35:43:@21.10]
  assign _GEN_11 = 5'hb == io_write_sel ? io_write_data : register_file_block_11; // @[regFile.scala 35:43:@21.10]
  assign _GEN_12 = 5'hc == io_write_sel ? io_write_data : register_file_block_12; // @[regFile.scala 35:43:@21.10]
  assign _GEN_13 = 5'hd == io_write_sel ? io_write_data : register_file_block_13; // @[regFile.scala 35:43:@21.10]
  assign _GEN_14 = 5'he == io_write_sel ? io_write_data : register_file_block_14; // @[regFile.scala 35:43:@21.10]
  assign _GEN_15 = 5'hf == io_write_sel ? io_write_data : register_file_block_15; // @[regFile.scala 35:43:@21.10]
  assign _GEN_16 = 5'h10 == io_write_sel ? io_write_data : register_file_block_16; // @[regFile.scala 35:43:@21.10]
  assign _GEN_17 = 5'h11 == io_write_sel ? io_write_data : register_file_block_17; // @[regFile.scala 35:43:@21.10]
  assign _GEN_18 = 5'h12 == io_write_sel ? io_write_data : register_file_block_18; // @[regFile.scala 35:43:@21.10]
  assign _GEN_19 = 5'h13 == io_write_sel ? io_write_data : register_file_block_19; // @[regFile.scala 35:43:@21.10]
  assign _GEN_20 = 5'h14 == io_write_sel ? io_write_data : register_file_block_20; // @[regFile.scala 35:43:@21.10]
  assign _GEN_21 = 5'h15 == io_write_sel ? io_write_data : register_file_block_21; // @[regFile.scala 35:43:@21.10]
  assign _GEN_22 = 5'h16 == io_write_sel ? io_write_data : register_file_block_22; // @[regFile.scala 35:43:@21.10]
  assign _GEN_23 = 5'h17 == io_write_sel ? io_write_data : register_file_block_23; // @[regFile.scala 35:43:@21.10]
  assign _GEN_24 = 5'h18 == io_write_sel ? io_write_data : register_file_block_24; // @[regFile.scala 35:43:@21.10]
  assign _GEN_25 = 5'h19 == io_write_sel ? io_write_data : register_file_block_25; // @[regFile.scala 35:43:@21.10]
  assign _GEN_26 = 5'h1a == io_write_sel ? io_write_data : register_file_block_26; // @[regFile.scala 35:43:@21.10]
  assign _GEN_27 = 5'h1b == io_write_sel ? io_write_data : register_file_block_27; // @[regFile.scala 35:43:@21.10]
  assign _GEN_28 = 5'h1c == io_write_sel ? io_write_data : register_file_block_28; // @[regFile.scala 35:43:@21.10]
  assign _GEN_29 = 5'h1d == io_write_sel ? io_write_data : register_file_block_29; // @[regFile.scala 35:43:@21.10]
  assign _GEN_30 = 5'h1e == io_write_sel ? io_write_data : register_file_block_30; // @[regFile.scala 35:43:@21.10]
  assign _GEN_31 = 5'h1f == io_write_sel ? io_write_data : register_file_block_31; // @[regFile.scala 35:43:@21.10]
  assign _GEN_32 = _T_68 ? _GEN_0 : 32'h0; // @[regFile.scala 34:53:@20.8]
  assign _GEN_33 = _T_68 ? _GEN_1 : register_file_block_1; // @[regFile.scala 34:53:@20.8]
  assign _GEN_34 = _T_68 ? _GEN_2 : register_file_block_2; // @[regFile.scala 34:53:@20.8]
  assign _GEN_35 = _T_68 ? _GEN_3 : register_file_block_3; // @[regFile.scala 34:53:@20.8]
  assign _GEN_36 = _T_68 ? _GEN_4 : register_file_block_4; // @[regFile.scala 34:53:@20.8]
  assign _GEN_37 = _T_68 ? _GEN_5 : register_file_block_5; // @[regFile.scala 34:53:@20.8]
  assign _GEN_38 = _T_68 ? _GEN_6 : register_file_block_6; // @[regFile.scala 34:53:@20.8]
  assign _GEN_39 = _T_68 ? _GEN_7 : register_file_block_7; // @[regFile.scala 34:53:@20.8]
  assign _GEN_40 = _T_68 ? _GEN_8 : register_file_block_8; // @[regFile.scala 34:53:@20.8]
  assign _GEN_41 = _T_68 ? _GEN_9 : register_file_block_9; // @[regFile.scala 34:53:@20.8]
  assign _GEN_42 = _T_68 ? _GEN_10 : register_file_block_10; // @[regFile.scala 34:53:@20.8]
  assign _GEN_43 = _T_68 ? _GEN_11 : register_file_block_11; // @[regFile.scala 34:53:@20.8]
  assign _GEN_44 = _T_68 ? _GEN_12 : register_file_block_12; // @[regFile.scala 34:53:@20.8]
  assign _GEN_45 = _T_68 ? _GEN_13 : register_file_block_13; // @[regFile.scala 34:53:@20.8]
  assign _GEN_46 = _T_68 ? _GEN_14 : register_file_block_14; // @[regFile.scala 34:53:@20.8]
  assign _GEN_47 = _T_68 ? _GEN_15 : register_file_block_15; // @[regFile.scala 34:53:@20.8]
  assign _GEN_48 = _T_68 ? _GEN_16 : register_file_block_16; // @[regFile.scala 34:53:@20.8]
  assign _GEN_49 = _T_68 ? _GEN_17 : register_file_block_17; // @[regFile.scala 34:53:@20.8]
  assign _GEN_50 = _T_68 ? _GEN_18 : register_file_block_18; // @[regFile.scala 34:53:@20.8]
  assign _GEN_51 = _T_68 ? _GEN_19 : register_file_block_19; // @[regFile.scala 34:53:@20.8]
  assign _GEN_52 = _T_68 ? _GEN_20 : register_file_block_20; // @[regFile.scala 34:53:@20.8]
  assign _GEN_53 = _T_68 ? _GEN_21 : register_file_block_21; // @[regFile.scala 34:53:@20.8]
  assign _GEN_54 = _T_68 ? _GEN_22 : register_file_block_22; // @[regFile.scala 34:53:@20.8]
  assign _GEN_55 = _T_68 ? _GEN_23 : register_file_block_23; // @[regFile.scala 34:53:@20.8]
  assign _GEN_56 = _T_68 ? _GEN_24 : register_file_block_24; // @[regFile.scala 34:53:@20.8]
  assign _GEN_57 = _T_68 ? _GEN_25 : register_file_block_25; // @[regFile.scala 34:53:@20.8]
  assign _GEN_58 = _T_68 ? _GEN_26 : register_file_block_26; // @[regFile.scala 34:53:@20.8]
  assign _GEN_59 = _T_68 ? _GEN_27 : register_file_block_27; // @[regFile.scala 34:53:@20.8]
  assign _GEN_60 = _T_68 ? _GEN_28 : register_file_block_28; // @[regFile.scala 34:53:@20.8]
  assign _GEN_61 = _T_68 ? _GEN_29 : register_file_block_29; // @[regFile.scala 34:53:@20.8]
  assign _GEN_62 = _T_68 ? _GEN_30 : register_file_block_30; // @[regFile.scala 34:53:@20.8]
  assign _GEN_63 = _T_68 ? _GEN_31 : register_file_block_31; // @[regFile.scala 34:53:@20.8]
  assign _GEN_64 = reset ? 32'h0 : _GEN_32; // @[regFile.scala 31:23:@13.6]
  assign _GEN_65 = reset ? register_file_block_1 : _GEN_33; // @[regFile.scala 31:23:@13.6]
  assign _GEN_66 = reset ? register_file_block_2 : _GEN_34; // @[regFile.scala 31:23:@13.6]
  assign _GEN_67 = reset ? register_file_block_3 : _GEN_35; // @[regFile.scala 31:23:@13.6]
  assign _GEN_68 = reset ? register_file_block_4 : _GEN_36; // @[regFile.scala 31:23:@13.6]
  assign _GEN_69 = reset ? register_file_block_5 : _GEN_37; // @[regFile.scala 31:23:@13.6]
  assign _GEN_70 = reset ? register_file_block_6 : _GEN_38; // @[regFile.scala 31:23:@13.6]
  assign _GEN_71 = reset ? register_file_block_7 : _GEN_39; // @[regFile.scala 31:23:@13.6]
  assign _GEN_72 = reset ? register_file_block_8 : _GEN_40; // @[regFile.scala 31:23:@13.6]
  assign _GEN_73 = reset ? register_file_block_9 : _GEN_41; // @[regFile.scala 31:23:@13.6]
  assign _GEN_74 = reset ? register_file_block_10 : _GEN_42; // @[regFile.scala 31:23:@13.6]
  assign _GEN_75 = reset ? register_file_block_11 : _GEN_43; // @[regFile.scala 31:23:@13.6]
  assign _GEN_76 = reset ? register_file_block_12 : _GEN_44; // @[regFile.scala 31:23:@13.6]
  assign _GEN_77 = reset ? register_file_block_13 : _GEN_45; // @[regFile.scala 31:23:@13.6]
  assign _GEN_78 = reset ? register_file_block_14 : _GEN_46; // @[regFile.scala 31:23:@13.6]
  assign _GEN_79 = reset ? register_file_block_15 : _GEN_47; // @[regFile.scala 31:23:@13.6]
  assign _GEN_80 = reset ? register_file_block_16 : _GEN_48; // @[regFile.scala 31:23:@13.6]
  assign _GEN_81 = reset ? register_file_block_17 : _GEN_49; // @[regFile.scala 31:23:@13.6]
  assign _GEN_82 = reset ? register_file_block_18 : _GEN_50; // @[regFile.scala 31:23:@13.6]
  assign _GEN_83 = reset ? register_file_block_19 : _GEN_51; // @[regFile.scala 31:23:@13.6]
  assign _GEN_84 = reset ? register_file_block_20 : _GEN_52; // @[regFile.scala 31:23:@13.6]
  assign _GEN_85 = reset ? register_file_block_21 : _GEN_53; // @[regFile.scala 31:23:@13.6]
  assign _GEN_86 = reset ? register_file_block_22 : _GEN_54; // @[regFile.scala 31:23:@13.6]
  assign _GEN_87 = reset ? register_file_block_23 : _GEN_55; // @[regFile.scala 31:23:@13.6]
  assign _GEN_88 = reset ? register_file_block_24 : _GEN_56; // @[regFile.scala 31:23:@13.6]
  assign _GEN_89 = reset ? register_file_block_25 : _GEN_57; // @[regFile.scala 31:23:@13.6]
  assign _GEN_90 = reset ? register_file_block_26 : _GEN_58; // @[regFile.scala 31:23:@13.6]
  assign _GEN_91 = reset ? register_file_block_27 : _GEN_59; // @[regFile.scala 31:23:@13.6]
  assign _GEN_92 = reset ? register_file_block_28 : _GEN_60; // @[regFile.scala 31:23:@13.6]
  assign _GEN_93 = reset ? register_file_block_29 : _GEN_61; // @[regFile.scala 31:23:@13.6]
  assign _GEN_94 = reset ? register_file_block_30 : _GEN_62; // @[regFile.scala 31:23:@13.6]
  assign _GEN_95 = reset ? register_file_block_31 : _GEN_63; // @[regFile.scala 31:23:@13.6]
  assign _GEN_129 = 5'h1 == io_read_sel1 ? register_file_block_1 : register_file_block_0; // @[regFile.scala 43:17:@28.4]
  assign _GEN_130 = 5'h2 == io_read_sel1 ? register_file_block_2 : _GEN_129; // @[regFile.scala 43:17:@28.4]
  assign _GEN_131 = 5'h3 == io_read_sel1 ? register_file_block_3 : _GEN_130; // @[regFile.scala 43:17:@28.4]
  assign _GEN_132 = 5'h4 == io_read_sel1 ? register_file_block_4 : _GEN_131; // @[regFile.scala 43:17:@28.4]
  assign _GEN_133 = 5'h5 == io_read_sel1 ? register_file_block_5 : _GEN_132; // @[regFile.scala 43:17:@28.4]
  assign _GEN_134 = 5'h6 == io_read_sel1 ? register_file_block_6 : _GEN_133; // @[regFile.scala 43:17:@28.4]
  assign _GEN_135 = 5'h7 == io_read_sel1 ? register_file_block_7 : _GEN_134; // @[regFile.scala 43:17:@28.4]
  assign _GEN_136 = 5'h8 == io_read_sel1 ? register_file_block_8 : _GEN_135; // @[regFile.scala 43:17:@28.4]
  assign _GEN_137 = 5'h9 == io_read_sel1 ? register_file_block_9 : _GEN_136; // @[regFile.scala 43:17:@28.4]
  assign _GEN_138 = 5'ha == io_read_sel1 ? register_file_block_10 : _GEN_137; // @[regFile.scala 43:17:@28.4]
  assign _GEN_139 = 5'hb == io_read_sel1 ? register_file_block_11 : _GEN_138; // @[regFile.scala 43:17:@28.4]
  assign _GEN_140 = 5'hc == io_read_sel1 ? register_file_block_12 : _GEN_139; // @[regFile.scala 43:17:@28.4]
  assign _GEN_141 = 5'hd == io_read_sel1 ? register_file_block_13 : _GEN_140; // @[regFile.scala 43:17:@28.4]
  assign _GEN_142 = 5'he == io_read_sel1 ? register_file_block_14 : _GEN_141; // @[regFile.scala 43:17:@28.4]
  assign _GEN_143 = 5'hf == io_read_sel1 ? register_file_block_15 : _GEN_142; // @[regFile.scala 43:17:@28.4]
  assign _GEN_144 = 5'h10 == io_read_sel1 ? register_file_block_16 : _GEN_143; // @[regFile.scala 43:17:@28.4]
  assign _GEN_145 = 5'h11 == io_read_sel1 ? register_file_block_17 : _GEN_144; // @[regFile.scala 43:17:@28.4]
  assign _GEN_146 = 5'h12 == io_read_sel1 ? register_file_block_18 : _GEN_145; // @[regFile.scala 43:17:@28.4]
  assign _GEN_147 = 5'h13 == io_read_sel1 ? register_file_block_19 : _GEN_146; // @[regFile.scala 43:17:@28.4]
  assign _GEN_148 = 5'h14 == io_read_sel1 ? register_file_block_20 : _GEN_147; // @[regFile.scala 43:17:@28.4]
  assign _GEN_149 = 5'h15 == io_read_sel1 ? register_file_block_21 : _GEN_148; // @[regFile.scala 43:17:@28.4]
  assign _GEN_150 = 5'h16 == io_read_sel1 ? register_file_block_22 : _GEN_149; // @[regFile.scala 43:17:@28.4]
  assign _GEN_151 = 5'h17 == io_read_sel1 ? register_file_block_23 : _GEN_150; // @[regFile.scala 43:17:@28.4]
  assign _GEN_152 = 5'h18 == io_read_sel1 ? register_file_block_24 : _GEN_151; // @[regFile.scala 43:17:@28.4]
  assign _GEN_153 = 5'h19 == io_read_sel1 ? register_file_block_25 : _GEN_152; // @[regFile.scala 43:17:@28.4]
  assign _GEN_154 = 5'h1a == io_read_sel1 ? register_file_block_26 : _GEN_153; // @[regFile.scala 43:17:@28.4]
  assign _GEN_155 = 5'h1b == io_read_sel1 ? register_file_block_27 : _GEN_154; // @[regFile.scala 43:17:@28.4]
  assign _GEN_156 = 5'h1c == io_read_sel1 ? register_file_block_28 : _GEN_155; // @[regFile.scala 43:17:@28.4]
  assign _GEN_157 = 5'h1d == io_read_sel1 ? register_file_block_29 : _GEN_156; // @[regFile.scala 43:17:@28.4]
  assign _GEN_158 = 5'h1e == io_read_sel1 ? register_file_block_30 : _GEN_157; // @[regFile.scala 43:17:@28.4]
  assign _GEN_161 = 5'h1 == io_read_sel2 ? register_file_block_1 : register_file_block_0; // @[regFile.scala 44:17:@29.4]
  assign _GEN_162 = 5'h2 == io_read_sel2 ? register_file_block_2 : _GEN_161; // @[regFile.scala 44:17:@29.4]
  assign _GEN_163 = 5'h3 == io_read_sel2 ? register_file_block_3 : _GEN_162; // @[regFile.scala 44:17:@29.4]
  assign _GEN_164 = 5'h4 == io_read_sel2 ? register_file_block_4 : _GEN_163; // @[regFile.scala 44:17:@29.4]
  assign _GEN_165 = 5'h5 == io_read_sel2 ? register_file_block_5 : _GEN_164; // @[regFile.scala 44:17:@29.4]
  assign _GEN_166 = 5'h6 == io_read_sel2 ? register_file_block_6 : _GEN_165; // @[regFile.scala 44:17:@29.4]
  assign _GEN_167 = 5'h7 == io_read_sel2 ? register_file_block_7 : _GEN_166; // @[regFile.scala 44:17:@29.4]
  assign _GEN_168 = 5'h8 == io_read_sel2 ? register_file_block_8 : _GEN_167; // @[regFile.scala 44:17:@29.4]
  assign _GEN_169 = 5'h9 == io_read_sel2 ? register_file_block_9 : _GEN_168; // @[regFile.scala 44:17:@29.4]
  assign _GEN_170 = 5'ha == io_read_sel2 ? register_file_block_10 : _GEN_169; // @[regFile.scala 44:17:@29.4]
  assign _GEN_171 = 5'hb == io_read_sel2 ? register_file_block_11 : _GEN_170; // @[regFile.scala 44:17:@29.4]
  assign _GEN_172 = 5'hc == io_read_sel2 ? register_file_block_12 : _GEN_171; // @[regFile.scala 44:17:@29.4]
  assign _GEN_173 = 5'hd == io_read_sel2 ? register_file_block_13 : _GEN_172; // @[regFile.scala 44:17:@29.4]
  assign _GEN_174 = 5'he == io_read_sel2 ? register_file_block_14 : _GEN_173; // @[regFile.scala 44:17:@29.4]
  assign _GEN_175 = 5'hf == io_read_sel2 ? register_file_block_15 : _GEN_174; // @[regFile.scala 44:17:@29.4]
  assign _GEN_176 = 5'h10 == io_read_sel2 ? register_file_block_16 : _GEN_175; // @[regFile.scala 44:17:@29.4]
  assign _GEN_177 = 5'h11 == io_read_sel2 ? register_file_block_17 : _GEN_176; // @[regFile.scala 44:17:@29.4]
  assign _GEN_178 = 5'h12 == io_read_sel2 ? register_file_block_18 : _GEN_177; // @[regFile.scala 44:17:@29.4]
  assign _GEN_179 = 5'h13 == io_read_sel2 ? register_file_block_19 : _GEN_178; // @[regFile.scala 44:17:@29.4]
  assign _GEN_180 = 5'h14 == io_read_sel2 ? register_file_block_20 : _GEN_179; // @[regFile.scala 44:17:@29.4]
  assign _GEN_181 = 5'h15 == io_read_sel2 ? register_file_block_21 : _GEN_180; // @[regFile.scala 44:17:@29.4]
  assign _GEN_182 = 5'h16 == io_read_sel2 ? register_file_block_22 : _GEN_181; // @[regFile.scala 44:17:@29.4]
  assign _GEN_183 = 5'h17 == io_read_sel2 ? register_file_block_23 : _GEN_182; // @[regFile.scala 44:17:@29.4]
  assign _GEN_184 = 5'h18 == io_read_sel2 ? register_file_block_24 : _GEN_183; // @[regFile.scala 44:17:@29.4]
  assign _GEN_185 = 5'h19 == io_read_sel2 ? register_file_block_25 : _GEN_184; // @[regFile.scala 44:17:@29.4]
  assign _GEN_186 = 5'h1a == io_read_sel2 ? register_file_block_26 : _GEN_185; // @[regFile.scala 44:17:@29.4]
  assign _GEN_187 = 5'h1b == io_read_sel2 ? register_file_block_27 : _GEN_186; // @[regFile.scala 44:17:@29.4]
  assign _GEN_188 = 5'h1c == io_read_sel2 ? register_file_block_28 : _GEN_187; // @[regFile.scala 44:17:@29.4]
  assign _GEN_189 = 5'h1d == io_read_sel2 ? register_file_block_29 : _GEN_188; // @[regFile.scala 44:17:@29.4]
  assign _GEN_190 = 5'h1e == io_read_sel2 ? register_file_block_30 : _GEN_189; // @[regFile.scala 44:17:@29.4]
  assign io_read_data1 = 5'h1f == io_read_sel1 ? register_file_block_31 : _GEN_158; // @[regFile.scala 43:17:@28.4]
  assign io_read_data2 = 5'h1f == io_read_sel2 ? register_file_block_31 : _GEN_190; // @[regFile.scala 44:17:@29.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  register_file_block_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  register_file_block_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  register_file_block_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  register_file_block_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  register_file_block_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  register_file_block_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  register_file_block_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  register_file_block_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  register_file_block_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  register_file_block_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  register_file_block_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  register_file_block_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  register_file_block_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  register_file_block_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  register_file_block_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  register_file_block_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  register_file_block_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  register_file_block_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  register_file_block_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  register_file_block_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  register_file_block_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  register_file_block_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  register_file_block_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  register_file_block_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  register_file_block_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  register_file_block_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  register_file_block_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  register_file_block_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  register_file_block_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  register_file_block_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  register_file_block_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  register_file_block_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_60) begin
      if (reset) begin
        register_file_block_0 <= 32'h0;
      end else begin
        if (_T_68) begin
          if (5'h0 == io_write_sel) begin
            register_file_block_0 <= io_write_data;
          end
        end else begin
          register_file_block_0 <= 32'h0;
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1 == io_write_sel) begin
            register_file_block_1 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h2 == io_write_sel) begin
            register_file_block_2 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h3 == io_write_sel) begin
            register_file_block_3 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h4 == io_write_sel) begin
            register_file_block_4 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h5 == io_write_sel) begin
            register_file_block_5 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h6 == io_write_sel) begin
            register_file_block_6 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h7 == io_write_sel) begin
            register_file_block_7 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h8 == io_write_sel) begin
            register_file_block_8 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h9 == io_write_sel) begin
            register_file_block_9 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'ha == io_write_sel) begin
            register_file_block_10 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'hb == io_write_sel) begin
            register_file_block_11 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'hc == io_write_sel) begin
            register_file_block_12 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'hd == io_write_sel) begin
            register_file_block_13 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'he == io_write_sel) begin
            register_file_block_14 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'hf == io_write_sel) begin
            register_file_block_15 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h10 == io_write_sel) begin
            register_file_block_16 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h11 == io_write_sel) begin
            register_file_block_17 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h12 == io_write_sel) begin
            register_file_block_18 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h13 == io_write_sel) begin
            register_file_block_19 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h14 == io_write_sel) begin
            register_file_block_20 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h15 == io_write_sel) begin
            register_file_block_21 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h16 == io_write_sel) begin
            register_file_block_22 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h17 == io_write_sel) begin
            register_file_block_23 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h18 == io_write_sel) begin
            register_file_block_24 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h19 == io_write_sel) begin
            register_file_block_25 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1a == io_write_sel) begin
            register_file_block_26 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1b == io_write_sel) begin
            register_file_block_27 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1c == io_write_sel) begin
            register_file_block_28 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1d == io_write_sel) begin
            register_file_block_29 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1e == io_write_sel) begin
            register_file_block_30 <= io_write_data;
          end
        end
      end
    end
    if (_T_60) begin
      if (!(reset)) begin
        if (_T_68) begin
          if (5'h1f == io_write_sel) begin
            register_file_block_31 <= io_write_data;
          end
        end
      end
    end
  end
endmodule
